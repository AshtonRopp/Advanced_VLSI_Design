`timescale 1ns/1ps

module Three_Parallel (
    input logic clk,
    input logic rst,
    input logic signed [15:0] din1,
    input logic signed [15:0] din2,
    input logic signed [15:0] din3,
    output logic signed [63:0] dout1,
    output logic signed [63:0] dout2,
    output logic signed [63:0] dout3
);

    localparam int TAPS = 102;

    // Buffers to store the most recent 102 samples
    logic signed [15:0] buffer0 [TAPS/3-1:0];
    logic signed [15:0] buffer1 [TAPS/3-1:0];
    logic signed [15:0] buffer2 [TAPS/3-1:0];
    
    // Coefficients for the FIR filter
    logic signed [31:0] H0 [TAPS/3-1:0];
    logic signed [31:0] H1 [TAPS/3-1:0];
    logic signed [31:0] H2 [TAPS/3-1:0];

    logic signed [31:0] coef [TAPS-1:0] = '{
            32'b11111111111110000101000100011100,
            32'b11111111111000110010100001001110,
            32'b11111111101101000000010001110011,
            32'b11111111010111011101110000111000,
            32'b11111110110101011110110010000100,
            32'b11111110000110010100100000001110,
            32'b11111101001100100110001111000010,
            32'b11111100001111001011001111010110,
            32'b11111011011001000010101110010000,
            32'b11111010110111110010101000110100,
            32'b11111010111000101110000110111000,
            32'b11111011100101000100011110011001,
            32'b11111100111110010111010100010101,
            32'b11111110111100000101010000001000,
            32'b00000001001011101110100110110101,
            32'b00000011010011110110001000001100,
            32'b00000100111001101000100110000110,
            32'b00000101100111111010111100110001,
            32'b00000101010101100010100111100101,
            32'b00000100001001000010111110000001,
            32'b00000010011000001101001000111111,
            32'b00000000100010111001101111101100,
            32'b11111111001010100000100110100001,
            32'b11111110101000000110001000011001,
            32'b11111111000100011111011111101110,
            32'b00000000010100111100110110111100,
            32'b00000001111101110111111000010001,
            32'b00000011011011001011111111100001,
            32'b00000100001100000000101100011010,
            32'b00000011111101111001110010001101,
            32'b00000010110011110110100011111110,
            32'b00000001000110010010100000101101,
            32'b11111111011011100111010000000100,
            32'b11111110011011010011001101101110,
            32'b11111110011111101100110010101111,
            32'b11111111101011011100101000111111,
            32'b00000001100110100010000111100001,
            32'b00000011100100101110100110111001,
            32'b00000100110011111011100110100011,
            32'b00000100101110000110100000111010,
            32'b00000011001000110110001101011100,
            32'b00000000011101000010001100100101,
            32'b11111101100011000100010101000111,
            32'b11111011100100000011000000011100,
            32'b11111011100011110001010101110010,
            32'b11111110001010001101000101110100,
            32'b00000011010011101001110010101011,
            32'b00001010001101001001100110000011,
            32'b00010001011110111100101000011100,
            32'b00010111100010100111010001011110,
            32'b00011010111110100000001110101110,
            32'b00011010111110100000001110101110,
            32'b00010111100010100111010001011110,
            32'b00010001011110111100101000011100,
            32'b00001010001101001001100110000011,
            32'b00000011010011101001110010101011,
            32'b11111110001010001101000101110100,
            32'b11111011100011110001010101110010,
            32'b11111011100100000011000000011100,
            32'b11111101100011000100010101000111,
            32'b00000000011101000010001100100101,
            32'b00000011001000110110001101011100,
            32'b00000100101110000110100000111010,
            32'b00000100110011111011100110100011,
            32'b00000011100100101110100110111001,
            32'b00000001100110100010000111100001,
            32'b11111111101011011100101000111111,
            32'b11111110011111101100110010101111,
            32'b11111110011011010011001101101110,
            32'b11111111011011100111010000000100,
            32'b00000001000110010010100000101101,
            32'b00000010110011110110100011111110,
            32'b00000011111101111001110010001101,
            32'b00000100001100000000101100011010,
            32'b00000011011011001011111111100001,
            32'b00000001111101110111111000010001,
            32'b00000000010100111100110110111100,
            32'b11111111000100011111011111101110,
            32'b11111110101000000110001000011001,
            32'b11111111001010100000100110100001,
            32'b00000000100010111001101111101100,
            32'b00000010011000001101001000111111,
            32'b00000100001001000010111110000001,
            32'b00000101010101100010100111100101,
            32'b00000101100111111010111100110001,
            32'b00000100111001101000100110000110,
            32'b00000011010011110110001000001100,
            32'b00000001001011101110100110110101,
            32'b11111110111100000101010000001000,
            32'b11111100111110010111010100010101,
            32'b11111011100101000100011110011001,
            32'b11111010111000101110000110111000,
            32'b11111010110111110010101000110100,
            32'b11111011011001000010101110010000,
            32'b11111100001111001011001111010110,
            32'b11111101001100100110001111000010,
            32'b11111110000110010100100000001110,
            32'b11111110110101011110110010000100,
            32'b11111111010111011101110000111000,
            32'b11111111101101000000010001110011,
            32'b11111111111000110010100001001110,
            32'b11111111111110000101000100011100
        };

    // Filter sums
    logic signed [63:0] sum_h0, sum_h1, sum_h2, sum_h01, sum_h12, sum_h012, sum_h2_reg, add_h1h2_min_h1_reg;
    logic signed [63:0] add_h01_min_h1, add_h12_min_h1, add_h012_min_add_h01_min_h1, add_h0_min_sum_h2_reg;

    // Assign adder outputs (excluding those attached to an output)
    assign add_h01_min_h1 = sum_h01 - sum_h1;
    assign add_h12_min_h1 = sum_h12 - sum_h1;
    assign add_h012_min_add_h01_min_h1 = sum_h012 - add_h01_min_h1;
    assign add_h0_min_sum_h2_reg = sum_h0 - sum_h2_reg;

    // Read coefficients from file
    always_comb begin
        for (int i = 0; 3*i < TAPS; i++) begin
            H0[i] = coef[3*i];
            
            if (3*i+1 < TAPS) begin
                H1[i] = coef[3*i+1];
            end
            if (3*i+2 < TAPS) begin
                H2[i] = coef[3*i+2];
            end
        end
    end

    // Process inputs
    always_ff @(posedge clk or posedge rst) begin
        if (rst) begin
            sum_h2_reg <= 0;
            add_h1h2_min_h1_reg <= 0;
            for (int i = 0; i <= TAPS/3-1; i++) begin
                buffer0[i] <= 0;
                buffer1[i] <= 0;
                buffer2[i] <= 0;
            end
        end
        else begin
            // Shift buffer and insert new input sample
            for (int i = TAPS/3-1; i > 0; i--) begin
                buffer0[i] <= buffer0[i - 1];
                buffer1[i] <= buffer1[i - 1];
                buffer2[i] <= buffer2[i - 1];
            end
            buffer0[0] <= din1;
            buffer1[0] <= din2;
            buffer2[0] <= din3;

            sum_h2_reg <= sum_h2;
            add_h1h2_min_h1_reg <= add_h12_min_h1;
        end
    end

    always_comb begin
        sum_h0 = 0;
        sum_h1 = 0;
        sum_h2 = 0;
        sum_h01 = 0;
        sum_h12 = 0;
        sum_h012 = 0;

        for (int i = 0; i <= TAPS/3-1; i++) begin
            sum_h0 += buffer0[i] * H0[i];
            sum_h1 += buffer1[i] * H1[i];
            sum_h2 += buffer2[i] * H2[i];

            sum_h01  += (buffer0[i] + buffer1[i])*(H0[i] + H1[i]);
            sum_h12  += (buffer1[i] + buffer2[i])*(H1[i] + H2[i]);
            sum_h012 += (buffer0[i] + buffer1[i] + buffer2[i])*(H0[i] + H1[i] + H2[i]);
        end
    end

    // Assign final outputs
    assign dout1 = (add_h0_min_sum_h2_reg + add_h1h2_min_h1_reg) >>> 31;
    assign dout2 = (add_h01_min_h1 - add_h0_min_sum_h2_reg) >>> 31;
    assign dout3 = (add_h012_min_add_h01_min_h1 - add_h12_min_h1) >>> 31;

endmodule
